
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);

-- GENERATED BY BC_MEM_PACKER
-- DATE: Mon Jun 06 17:39:44 2016

	signal mem : ram_t := (
		-- Tile Matrix
		0 => x"00000001",
		1 => x"00000000",
		2 => x"00000001",
		3 => x"00000000",
		4 => x"00000001",
		5 => x"00000000",
		6 => x"00000001",
		7 => x"00000000",
		8 => x"00000001",
		9 => x"00000000",
		10 => x"00000001",
		11 => x"00000000",
		12 => x"00000001",
		13 => x"00000000",
		14 => x"00000001",
		15 => x"00000000",
		16 => x"00000001",
		17 => x"00000000",
		18 => x"00000001",
		19 => x"00000000",
		20 => x"00000001",
		21 => x"00000000",
		22 => x"00000001",
		23 => x"00000000",
		24 => x"00000001",
		25 => x"00000000", -----------
		26 => x"00000000",
		27 => x"00000000",
		28 => x"00000000",
		29 => x"00000000",
		30 => x"00000001",
		31 => x"00000000",
		32 => x"00000001",
		33 => x"00000000",
		34 => x"00000001",
		35 => x"00000000",
		36 => x"00000001",
		37 => x"00000000",
		38 => x"00000001",
		39 => x"00000000",
		40 => x"00000001",
		41 => x"00000000",
		42 => x"00000001",
		43 => x"00000000",
		44 => x"00000001",
		45 => x"00000000",
		46 => x"00000001",
		47 => x"00000000",
		48 => x"00000001",
		49 => x"00000000",
		50 => x"00000001",
		51 => x"00000000",
		52 => x"00000001",
		53 => x"00000000",
		54 => x"00000001",
		55 => x"00000000",
		56 => x"00000000",
		57 => x"00000000",
		58 => x"00000000",
		59 => x"00000000",
		60 => x"00000001",
		61 => x"00000000",
		62 => x"00000001",
		63 => x"00000000",
		64 => x"00000001",
		65 => x"00000000",
		66 => x"00000001",
		67 => x"00000000",
		68 => x"00000001",
		69 => x"00000000",
		70 => x"00000001",
		71 => x"00000000",
		72 => x"00000001",
		73 => x"00000000",
		74 => x"00000001",
		75 => x"00000000",
		76 => x"00000001",
		77 => x"00000000",
		78 => x"00000001",
		79 => x"00000000",
		80 => x"00000001",
		81 => x"00000000",
		82 => x"00000001",
		83 => x"00000000",
		84 => x"00000001",
		85 => x"00000000",
		86 => x"00000000",
		87 => x"00000000",
		88 => x"00000000",
		89 => x"00000000",
		90 => x"00000001",
		91 => x"00000000",
		92 => x"00000001",
		93 => x"00000000",
		94 => x"00000001",
		95 => x"00000000",
		96 => x"00000102", -----
		97 => x"00000000",
		98 => x"00000102",
		99 => x"00000000",
		100 => x"00000102",
		101 => x"00000000",
		102 => x"00000102",
		103 => x"00000000",
		104 => x"00000102",
		105 => x"00000000",
		106 => x"00000102",
		107 => x"00000000",
		108 => x"00000102",
		109 => x"00000000",
		110 => x"00000001",
		111 => x"00000000",
		112 => x"00000001",
		113 => x"00000000",
		114 => x"00000001",
		115 => x"00000000",
		116 => x"00000000",
		117 => x"00000000",
		118 => x"00000000",
		119 => x"00000000",
		120 => x"00000001",
		121 => x"00000000",
		122 => x"00000001",
		123 => x"00000000",
		124 => x"00000001",
		125 => x"00000000",
		126 => x"00000102",
		127 => x"00000000",
		128 => x"00000102",
		129 => x"00000000",
		130 => x"00000102",
		131 => x"00000000",
		132 => x"00000102",
		133 => x"00000000",
		134 => x"00000102",
		135 => x"00000000",
		136 => x"00000102",
		137 => x"00000000",
		138 => x"00000102",
		139 => x"00000000",
		140 => x"00000001",
		141 => x"00000000",
		142 => x"00000001",
		143 => x"00000000",
		144 => x"00000001",
		145 => x"00000000",
		146 => x"00000000",
		147 => x"00000000",
		148 => x"00000000",
		149 => x"00000000",
		150 => x"00000001",
		151 => x"00000000",
		152 => x"00000001",
		153 => x"00000000",
		154 => x"00000001",
		155 => x"00000000",
		156 => x"00000102",
		157 => x"00000000",
		158 => x"00000102",
		159 => x"00000000",
		160 => x"00000102",
		161 => x"00000000",
		162 => x"00000102",
		163 => x"00000000",
		164 => x"00000102",
		165 => x"00000000",
		166 => x"00000102",
		167 => x"00000000",
		168 => x"00000102",
		169 => x"00000000",
		170 => x"00000001",
		171 => x"00000000",
		172 => x"00000001",
		173 => x"00000000",
		174 => x"00000001",
		175 => x"00000000",
		176 => x"00000000",
		177 => x"00000000",
		178 => x"00000000",
		179 => x"00000000",
		180 => x"00000001",
		181 => x"00000000",
		182 => x"00000001",
		183 => x"00000000",
		184 => x"00000001",
		185 => x"00000000",
		186 => x"00000102",
		187 => x"00000000",
		188 => x"00000102",
		189 => x"00000000",
		190 => x"00000102",
		191 => x"00000000",
		192 => x"00000102",
		193 => x"00000000",
		194 => x"00000102",
		195 => x"00000000",
		196 => x"00000102",
		197 => x"00000000",
		198 => x"00000102",
		199 => x"00000000",
		200 => x"00000001",
		201 => x"00000000",
		202 => x"00000001",
		203 => x"00000000",
		204 => x"00000001",
		205 => x"00000000",
		206 => x"00000000",
		207 => x"00000000",
		208 => x"00000000",
		209 => x"00000000",
		210 => x"00000001",
		211 => x"00000000",
		212 => x"00000001",
		213 => x"00000000",
		214 => x"00000001",
		215 => x"00000000",
		216 => x"00000102",
		217 => x"00000000",
		218 => x"00000102",
		219 => x"00000000",
		220 => x"00000102",
		221 => x"00000000",
		222 => x"00000102",
		223 => x"00000000",
		224 => x"00000102",
		225 => x"00000000",
		226 => x"00000102",
		227 => x"00000000",
		228 => x"00000102",
		229 => x"00000000",
		230 => x"00000001",
		231 => x"00000000",
		232 => x"00000001",
		233 => x"00000000",
		234 => x"00000001",
		235 => x"00000000",
		236 => x"00000000",
		237 => x"00000000",
		238 => x"00000000",
		239 => x"00000000",
		240 => x"00000001",
		241 => x"00000000",
		242 => x"00000001",
		243 => x"00000000",
		244 => x"00000001",
		245 => x"00000000",
		246 => x"00000001",
		247 => x"00000000",
		248 => x"00000001",
		249 => x"00000000",
		250 => x"00000001",
		251 => x"00000000",
		252 => x"00000001",
		253 => x"00000000",
		254 => x"00000001",
		255 => x"00000000",
		256 => x"00000001",
		257 => x"00000000",
		258 => x"00000001",
		259 => x"00000000",
		260 => x"00000001",
		261 => x"00000000",
		262 => x"00000001",
		263 => x"00000000",
		264 => x"00000001",
		265 => x"00000000",
		266 => x"00000000",
		267 => x"00000000",
		268 => x"00000000",
		269 => x"00000000",
		270 => x"00000001",
		271 => x"00000000",
		272 => x"00000001",
		273 => x"00000000",
		274 => x"00000001",
		275 => x"00000000",
		276 => x"00000202",
		277 => x"00000000",
		278 => x"00000202",
		279 => x"00000000",
		280 => x"00000202",
		281 => x"00000000",
		282 => x"00000202",
		283 => x"00000000",
		284 => x"00000202",
		285 => x"00000000",
		286 => x"00000202",
		287 => x"00000000",
		288 => x"00000202",
		289 => x"00000000",
		290 => x"00000001",
		291 => x"00000000",
		292 => x"00000001",
		293 => x"00000000",
		294 => x"00000001",
		295 => x"00000000",
		296 => x"00000000",
		297 => x"00000000",
		298 => x"00000000",
		299 => x"00000000",
		300 => x"00000001",
		301 => x"00000000",
		302 => x"00000001",
		303 => x"00000000",
		304 => x"00000001",
		305 => x"00000000",
		306 => x"00000202",
		307 => x"00000000",
		308 => x"00020303",
		309 => x"00000000",
		310 => x"00020303",
		311 => x"00000000",
		312 => x"00020303",
		313 => x"00000000",
		314 => x"00020303",
		315 => x"00000000",
		316 => x"00020303",
		317 => x"00000000",
		318 => x"00020303",
		319 => x"00000000",
		320 => x"00000302",
		321 => x"00000000",
		322 => x"00000302",
		323 => x"00000000",
		324 => x"00000302",
		325 => x"00000000",
		326 => x"00000301",
		327 => x"00000000",
		328 => x"00000301",
		329 => x"00000000",
		330 => x"00000001",
		331 => x"00000000",
		332 => x"00000001",
		333 => x"00000000",
		334 => x"00000001",
		335 => x"00000000",
		336 => x"00000202",
		337 => x"00000000",
		338 => x"00020303",
		339 => x"00000000",
		340 => x"00020303",
		341 => x"00000000",
		342 => x"00020303",
		343 => x"00000000",
		344 => x"00020303",
		345 => x"00000000",
		346 => x"00020303",
		347 => x"00000000",
		348 => x"00020303",
		349 => x"00000000",
		350 => x"00000302",
		351 => x"00000000",
		352 => x"00000302",
		353 => x"00000000",
		354 => x"00000302",
		355 => x"00000000",
		356 => x"00000301",
		357 => x"00000000",
		358 => x"00000301",
		359 => x"00000000",
		360 => x"00000001",
		361 => x"00000000",
		362 => x"00000001",
		363 => x"00000000",
		364 => x"00000001",
		365 => x"00000000",
		366 => x"00000202",
		367 => x"00000000",
		368 => x"00020303",
		369 => x"00000000",
		370 => x"00020303",
		371 => x"00000000",
		372 => x"02030404",
		373 => x"00000000",
		374 => x"02030404",
		375 => x"00000000",
		376 => x"02030404",
		377 => x"00000000",
		378 => x"02030404",
		379 => x"00000000",
		380 => x"00030403",
		381 => x"00000000",
		382 => x"00030403",
		383 => x"00000000",
		384 => x"00030403",
		385 => x"00000000",
		386 => x"00000301",
		387 => x"00000000",
		388 => x"00000301",
		389 => x"00000000",
		390 => x"00000001",
		391 => x"00000000",
		392 => x"00000001",
		393 => x"00000000",
		394 => x"00000001",
		395 => x"00000000",
		396 => x"00000202",
		397 => x"00000000",
		398 => x"00020303",
		399 => x"00000000",
		400 => x"00020303",
		401 => x"00000000",
		402 => x"02030404",
		403 => x"00000000",
		404 => x"02030404",   ----------------------------------------------------
		405 => x"00000000",
		406 => x"02030404",
		407 => x"00000000",
		408 => x"02030404",
		409 => x"00000000",
		410 => x"00030403",
		411 => x"00000000",
		412 => x"00030403",
		413 => x"00000000",
		414 => x"00030403",
		415 => x"00000000",
		416 => x"00000301",
		417 => x"00000000",
		418 => x"00000301",
		419 => x"00000000",
		420 => x"00000001",
		421 => x"00000000",
		422 => x"00000001",
		423 => x"00000000",
		424 => x"00000001",
		425 => x"00000000",
		426 => x"00000202",
		427 => x"00000000",
		428 => x"00020303",
		429 => x"00000000",
		430 => x"00020303",
		431 => x"00000000",
		432 => x"02030404",
		433 => x"00000000",
		434 => x"02030404",
		435 => x"00000000",
		436 => x"02030404",
		437 => x"00000000",
		438 => x"02030404",
		439 => x"00000000",
		440 => x"00030403",
		441 => x"00000000",
		442 => x"00030403",
		443 => x"00000000",
		444 => x"00030403",
		445 => x"00000000",
		446 => x"00000301",
		447 => x"00000000",
		448 => x"00000301",
		449 => x"00000000",
		450 => x"00000001",
		451 => x"00000000",
		452 => x"00000001",
		453 => x"00000000",
		454 => x"00000001",
		455 => x"00000000",
		456 => x"00000001",
		457 => x"00000000",
		458 => x"00000302",
		459 => x"00000000",
		460 => x"00000302",
		461 => x"00000000",
		462 => x"00030403",
		463 => x"00000000",
		464 => x"00030403",
		465 => x"00000000",
		466 => x"00030403",
		467 => x"00000000",
		468 => x"00030403",
		469 => x"00000000",
		470 => x"00030403",
		471 => x"00000000",
		472 => x"00030403",
		473 => x"00000000",
		474 => x"00030403",
		475 => x"00000000",
		476 => x"00000301",
		477 => x"00000000",
		478 => x"00000301",
		479 => x"00000000",
		480 => x"00000000",
		481 => x"00000000",
		482 => x"00000000",
		483 => x"00000000",
		484 => x"00000000",
		485 => x"00000000",
		486 => x"00000000",
		487 => x"00000000",
		488 => x"00000301",
		489 => x"00000000",
		490 => x"00000301",
		491 => x"00000000",
		492 => x"00030402",
		493 => x"00000000",
		494 => x"00030402",
		495 => x"00000000",
		496 => x"00030402",
		497 => x"00000000",
		498 => x"00030402",
		499 => x"00000000",
		500 => x"00030402",
		501 => x"00000000",
		502 => x"00030402",
		503 => x"00000000",
		504 => x"00030402",
		505 => x"00000000",
		506 => x"00000301",
		507 => x"00000000",
		508 => x"00000301",
		509 => x"00000000",
		510 => x"00000000",
		511 => x"00000000",
		512 => x"00000000",
		513 => x"00000000",
		514 => x"00000000",
		515 => x"00000000",
		516 => x"00000000",
		517 => x"00000000",
		518 => x"00000301",
		519 => x"00000000",
		520 => x"00000301",
		521 => x"00000000",
		522 => x"00030402",
		523 => x"00000000",
		524 => x"00030402",
		525 => x"00000000",
		526 => x"00030402",
		527 => x"00000000",
		528 => x"00030402",
		529 => x"00000000",
		530 => x"00030402",
		531 => x"00000000",
		532 => x"00030402",
		533 => x"00000000",
		534 => x"00030402",
		535 => x"00000000",
		536 => x"00000301",
		537 => x"00000000",
		538 => x"00000301",
		539 => x"00000000",
		540 => x"00000000",
		541 => x"00000000",
		542 => x"00000000",
		543 => x"00000000",
		544 => x"00000000",
		545 => x"00000000",
		546 => x"00000000",
		547 => x"00000000",
		548 => x"00000301",
		549 => x"00000000",
		550 => x"00000301",
		551 => x"00000000",
		552 => x"00030402",
		553 => x"00000000",
		554 => x"00030402",
		555 => x"00000000",
		556 => x"00030402",
		557 => x"00000000",
		558 => x"00030402",
		559 => x"00000000",
		560 => x"00030402",
		561 => x"00000000",
		562 => x"00030402",
		563 => x"00000000",
		564 => x"00030402",
		565 => x"00000000",
		566 => x"00000301",
		567 => x"00000000",
		568 => x"00000301",
		569 => x"00000000",
		570 => x"00000000",
		571 => x"00000000",
		572 => x"00000000",
		573 => x"00000000",
		574 => x"00000000",
		575 => x"00000000",
		576 => x"00000000",
		577 => x"00000000",
		578 => x"00000301",
		579 => x"00000000",
		580 => x"00000301",
		581 => x"00000000",
		582 => x"00000301",
		583 => x"00000000",
		584 => x"00000301",
		585 => x"00000000",
		586 => x"00000301",
		587 => x"00000000",
		588 => x"00000301",
		589 => x"00000000",
		590 => x"00000301",
		591 => x"00000000",
		592 => x"00000301",
		593 => x"00000000",
		594 => x"00000301",
		595 => x"00000000",
		596 => x"00000301",
		597 => x"00000000",
		598 => x"00000301",
		599 => x"00000000",
		-- Draw list
		600 => x"00000000",
		601 => x"019001f4",
		602 => x"00640064",
		603 => x"00c80096",
		604 => x"0064012c",
		605 => x"00c80096",
		606 => x"0096015e",
		607 => x"012c012c",
		608 => x"00c80190",
		609 => x"00c800c8",
		610 => x"00000000",
		611 => x"00000000",
		612 => x"00000000",
		613 => x"00000000",
		614 => x"00000000",
		615 => x"00000000",
		616 => x"00000000",
		617 => x"00000000",
		618 => x"00000000",
		619 => x"00000000",
		620 => x"00000000",
		621 => x"00000000",
		622 => x"00000000",
		623 => x"00000000",
		624 => x"00000000",
		625 => x"00000000",
		626 => x"00000000",
		627 => x"00000000",
		628 => x"00000000",
		629 => x"00000000",
		630 => x"00000000",
		631 => x"00000000",
		632 => x"00000000",
		633 => x"00000000",
		634 => x"00000000",
		635 => x"00000000",
		636 => x"00000000",
		637 => x"00000000",
		638 => x"00000000",
		639 => x"00000000",
		640 => x"00000000",
		641 => x"00000000",
		642 => x"00000000",
		643 => x"00000000",
		644 => x"00000000",
		645 => x"00000000",
		646 => x"00000000",
		647 => x"00000000",
		648 => x"00000000",
		649 => x"00000000",
		650 => x"00000000",
		651 => x"00000000",
		652 => x"00000000",
		653 => x"00000000",
		654 => x"00000000",
		655 => x"00000000",
		656 => x"00000000",
		657 => x"00000000",
		658 => x"00000000",
		659 => x"00000000",
		660 => x"00000000",
		661 => x"00000000",
		662 => x"00000000",
		663 => x"00000000",
		664 => x"00000000",
		665 => x"00000000",
		666 => x"00000000",
		667 => x"00000000",
		668 => x"00000000",
		669 => x"00000000",
		670 => x"00000000",
		671 => x"00000000",
		672 => x"00000000",
		673 => x"00000000",
		674 => x"00000000",
		675 => x"00000000",
		676 => x"00000000",
		677 => x"00000000",
		678 => x"00000000",
		679 => x"00000000",
		680 => x"00000000",
		681 => x"00000000",
		682 => x"00000000",
		683 => x"00000000",
		684 => x"00000000",
		685 => x"00000000",
		686 => x"00000000",
		687 => x"00000000",
		688 => x"00000000",
		689 => x"00000000",
		690 => x"00000000",
		691 => x"00000000",
		692 => x"00000000",
		693 => x"00000000",
		694 => x"00000000",
		695 => x"00000000",
		696 => x"00000000",
		697 => x"00000000",
		698 => x"00000000",
		699 => x"00000000",
		700 => x"00000000",
		701 => x"00000000",
		702 => x"00000000",
		703 => x"00000000",
		704 => x"00000000",
		705 => x"00000000",
		706 => x"00000000",
		707 => x"00000000",
		708 => x"00000000",
		709 => x"00000000",
		710 => x"00000000",
		711 => x"00000000",
		712 => x"00000000",
		713 => x"00000000",
		714 => x"00000000",
		715 => x"00000000",
		716 => x"00000000",
		717 => x"00000000",
		718 => x"00000000",
		719 => x"00000000",
		720 => x"00000000",
		721 => x"00000000",
		722 => x"00000000",
		723 => x"00000000",
		724 => x"00000000",
		725 => x"00000000",
		726 => x"00000000",
		727 => x"00000000",
		728 => x"00000000",
		729 => x"00000000",
		730 => x"00000000",
		731 => x"00000000",
		732 => x"00000000",
		733 => x"00000000",
		734 => x"00000000",
		735 => x"00000000",
		736 => x"00000000",
		737 => x"00000000",
		738 => x"00000000",
		739 => x"00000000",
		740 => x"00000000",
		741 => x"00000000",
		742 => x"00000000",
		743 => x"00000000",
		744 => x"00000000",
		745 => x"00000000",
		746 => x"00000000",
		747 => x"00000000",
		748 => x"00000000",
		749 => x"00000000",
		750 => x"00000000",
		751 => x"00000000",
		752 => x"00000000",
		753 => x"00000000",
		754 => x"00000000",
		755 => x"00000000",
		756 => x"00000000",
		757 => x"00000000",
		758 => x"00000000",
		759 => x"00000000",
		760 => x"00000000",
		761 => x"00000000",
		762 => x"00000000",
		763 => x"00000000",
		764 => x"00000000",
		765 => x"00000000",
		766 => x"00000000",
		767 => x"00000000",
		768 => x"00000000",
		769 => x"00000000",
		770 => x"00000000",
		771 => x"00000000",
		772 => x"00000000",
		773 => x"00000000",
		774 => x"00000000",
		775 => x"00000000",
		776 => x"00000000",
		777 => x"00000000",
		778 => x"00000000",
		779 => x"00000000",
		780 => x"00000000",
		781 => x"00000000",
		782 => x"00000000",
		783 => x"00000000",
		784 => x"00000000",
		785 => x"00000000",
		786 => x"00000000",
		787 => x"00000000",
		788 => x"00000000",
		789 => x"00000000",
		790 => x"00000000",
		791 => x"00000000",
		792 => x"00000000",
		793 => x"00000000",
		794 => x"00000000",
		795 => x"00000000",
		796 => x"00000000",
		797 => x"00000000",
		798 => x"00000000",
		799 => x"00000000",
		800 => x"00000000",
		801 => x"00000000",
		802 => x"00000000",
		803 => x"00000000",
		804 => x"00000000",
		805 => x"00000000",
		806 => x"00000000",
		807 => x"00000000",
		808 => x"00000000",
		809 => x"00000000",
		810 => x"00000000",
		811 => x"00000000",
		812 => x"00000000",
		813 => x"00000000",
		814 => x"00000000",
		815 => x"00000000",
		816 => x"00000000",
		817 => x"00000000",
		818 => x"00000000",
		819 => x"00000000",
		820 => x"00000000",
		821 => x"00000000",
		822 => x"00000000",
		823 => x"00000000",
		824 => x"00000000",
		825 => x"00000000",
		826 => x"00000000",
		827 => x"00000000",
		828 => x"00000000",
		829 => x"00000000",
		830 => x"00000000",
		831 => x"00000000",
		832 => x"00000000",
		833 => x"00000000",
		834 => x"00000000",
		835 => x"00000000",
		836 => x"00000000",
		837 => x"00000000",
		838 => x"00000000",
		839 => x"00000000",
		840 => x"00000000",
		841 => x"00000000",
		842 => x"00000000",
		843 => x"00000000",
		844 => x"00000000",
		845 => x"00000000",
		846 => x"00000000",
		847 => x"00000000",
		848 => x"00000000",
		849 => x"00000000",
		850 => x"00000000",
		851 => x"00000000",
		852 => x"00000000",
		853 => x"00000000",
		854 => x"00000000",
		855 => x"00000000",
		856 => x"00000000",
		857 => x"00000000",
		858 => x"00000000",
		859 => x"00000000",
		860 => x"00000000",
		861 => x"00000000",
		862 => x"00000000",
		863 => x"00000000",
		864 => x"00000000",
		865 => x"00000000",
		866 => x"00000000",
		867 => x"00000000",
		868 => x"00000000",
		869 => x"00000000",
		870 => x"00000000",
		871 => x"00000000",
		872 => x"00000000",
		873 => x"00000000",
		874 => x"00000000",
		875 => x"00000000",
		876 => x"00000000",
		877 => x"00000000",
		878 => x"00000000",
		879 => x"00000000",
		880 => x"00000000",
		881 => x"00000000",
		882 => x"00000000",
		883 => x"00000000",
		884 => x"00000000",
		885 => x"00000000",
		886 => x"00000000",
		887 => x"00000000",
		888 => x"00000000",
		889 => x"00000000",
		890 => x"00000000",
		891 => x"00000000",
		892 => x"00000000",
		893 => x"00000000",
		894 => x"00000000",
		895 => x"00000000",
		896 => x"00000000",
		897 => x"00000000",
		898 => x"00000000",
		899 => x"00000000",
		900 => x"00000000",
		901 => x"00000000",
		902 => x"00000000",
		903 => x"00000000",
		904 => x"00000000",
		905 => x"00000000",
		906 => x"00000000",
		907 => x"00000000",
		908 => x"00000000",
		909 => x"00000000",
		910 => x"00000000",
		911 => x"00000000",
		912 => x"00000000",
		913 => x"00000000",
		914 => x"00000000",
		915 => x"00000000",
		916 => x"00000000",
		917 => x"00000000",
		918 => x"00000000",
		919 => x"00000000",
		920 => x"00000000",
		921 => x"00000000",
		922 => x"00000000",
		923 => x"00000000",
		924 => x"00000000",
		925 => x"00000000",
		926 => x"00000000",
		927 => x"00000000",
		928 => x"00000000",
		929 => x"00000000",
		930 => x"00000000",
		931 => x"00000000",
		932 => x"00000000",
		933 => x"00000000",
		934 => x"00000000",
		935 => x"00000000",
		936 => x"00000000",
		937 => x"00000000",
		938 => x"00000000",
		939 => x"00000000",
		940 => x"00000000",
		941 => x"00000000",
		942 => x"00000000",
		943 => x"00000000",
		944 => x"00000000",
		945 => x"00000000",
		946 => x"00000000",
		947 => x"00000000",
		948 => x"00000000",
		949 => x"00000000",
		950 => x"00000000",
		951 => x"00000000",
		952 => x"00000000",
		953 => x"00000000",
		954 => x"00000000",
		955 => x"00000000",
		956 => x"00000000",
		957 => x"00000000",
		958 => x"00000000",
		959 => x"00000000",
		960 => x"00000000",
		961 => x"00000000",
		962 => x"00000000",
		963 => x"00000000",
		964 => x"00000000",
		965 => x"00000000",
		966 => x"00000000",
		967 => x"00000000",
		968 => x"00000000",
		969 => x"00000000",
		970 => x"00000000",
		971 => x"00000000",
		972 => x"00000000",
		973 => x"00000000",
		974 => x"00000000",
		975 => x"00000000",
		976 => x"00000000",
		977 => x"00000000",
		978 => x"00000000",
		979 => x"00000000",
		980 => x"00000000",
		981 => x"00000000",
		982 => x"00000000",
		983 => x"00000000",
		984 => x"00000000",
		985 => x"00000000",
		986 => x"00000000",
		987 => x"00000000",
		988 => x"00000000",
		989 => x"00000000",
		990 => x"00000000",
		991 => x"00000000",
		992 => x"00000000",
		993 => x"00000000",
		994 => x"00000000",
		995 => x"00000000",
		996 => x"00000000",
		997 => x"00000000",
		998 => x"00000000",
		999 => x"00000000",
		1000 => x"00000000",
		1001 => x"00000000",
		1002 => x"00000000",
		1003 => x"00000000",
		1004 => x"00000000",
		1005 => x"00000000",
		1006 => x"00000000",
		1007 => x"00000000",
		1008 => x"00000000",
		1009 => x"00000000",
		1010 => x"00000000",
		1011 => x"00000000",
		1012 => x"00000000",
		1013 => x"00000000",
		1014 => x"00000000",
		1015 => x"00000000",
		1016 => x"00000000",
		1017 => x"00000000",
		1018 => x"00000000",
		1019 => x"00000000",
		1020 => x"00000000",
		1021 => x"00000000",
		1022 => x"00000000",
		1023 => x"00000000",
		1024 => x"00000000",
		1025 => x"00000000",
		1026 => x"00000000",
		1027 => x"00000000",
		1028 => x"00000000",
		1029 => x"00000000",
		1030 => x"00000000",
		1031 => x"00000000",
		1032 => x"00000000",
		1033 => x"00000000",
		1034 => x"00000000",
		1035 => x"00000000",
		1036 => x"00000000",
		1037 => x"00000000",
		1038 => x"00000000",
		1039 => x"00000000",
		1040 => x"00000000",
		1041 => x"00000000",
		1042 => x"00000000",
		1043 => x"00000000",
		1044 => x"00000000",
		1045 => x"00000000",
		1046 => x"00000000",
		1047 => x"00000000",
		1048 => x"00000000",
		1049 => x"00000000",
		1050 => x"00000000",
		1051 => x"00000000",
		1052 => x"00000000",
		1053 => x"00000000",
		1054 => x"00000000",
		1055 => x"00000000",
		1056 => x"00000000",
		1057 => x"00000000",
		1058 => x"00000000",
		1059 => x"00000000",
		1060 => x"00000000",
		1061 => x"00000000",
		1062 => x"00000000",
		1063 => x"00000000",
		1064 => x"00000000",
		1065 => x"00000000",
		1066 => x"00000000",
		1067 => x"00000000",
		1068 => x"00000000",
		1069 => x"00000000",
		1070 => x"00000000",
		1071 => x"00000000",
		1072 => x"00000000",
		1073 => x"00000000",
		1074 => x"00000000",
		1075 => x"00000000",
		1076 => x"00000000",
		1077 => x"00000000",
		1078 => x"00000000",
		1079 => x"00000000",
		1080 => x"00000000",
		1081 => x"00000000",
		1082 => x"00000000",
		1083 => x"00000000",
		1084 => x"00000000",
		1085 => x"00000000",
		1086 => x"00000000",
		1087 => x"00000000",
		1088 => x"00000000",
		1089 => x"00000000",
		1090 => x"00000000",
		1091 => x"00000000",
		1092 => x"00000000",
		1093 => x"00000000",
		1094 => x"00000000",
		1095 => x"00000000",
		1096 => x"00000000",
		1097 => x"00000000",
		1098 => x"00000000",
		1099 => x"00000000",
		1100 => x"00000000",
		1101 => x"00000000",
		1102 => x"00000000",
		1103 => x"00000000",
		1104 => x"00000000",
		1105 => x"00000000",
		1106 => x"00000000",
		1107 => x"00000000",
		1108 => x"00000000",
		1109 => x"00000000",
		1110 => x"00000000",
		1111 => x"00000000",
		1112 => x"ff0000ff",
		1113 => x"ff8080ff",
		1114 => x"ff8080ff",
		1115 => x"80ff0000",
		1116 => x"ffff8080",
		1117 => x"00000000",
		1118 => x"00000000",
		1119 => x"00000000",
		1120 => x"00000000",
		1121 => x"00000000",
		1122 => x"00000000",
		1123 => x"00000000",
		1124 => x"00000000",
		1125 => x"00000000",
		1126 => x"00000000",
		1127 => x"00000000",
		1128 => x"00000000",
		1129 => x"00000000",
		1130 => x"00000000",
		1131 => x"00000000",
		1132 => x"00000000",
		1133 => x"00000000",
		1134 => x"00000000",
		1135 => x"00000000",
		1136 => x"00000000",
		1137 => x"00000000",
		1138 => x"00000000",
		1139 => x"00000000",
		1140 => x"00000000",
		1141 => x"00000000",
		1142 => x"00000000",
		1143 => x"00000000",
		1144 => x"00000000",
		1145 => x"00000000",
		1146 => x"00000000",
		1147 => x"00000000",
		1148 => x"00000000",
		1149 => x"00000000",
		1150 => x"00000000",
		1151 => x"00000000",
		1152 => x"00000000",
		1153 => x"00000000",
		1154 => x"00000000",
		1155 => x"00000000",
		1156 => x"00000000",
		1157 => x"00000000",
		1158 => x"00000000",
		1159 => x"00000000",
		1160 => x"00000000",
		1161 => x"00000000",
		1162 => x"00000000",
		1163 => x"00000000",
		1164 => x"00000000",
		1165 => x"00000000",
		1166 => x"00000000",
		1167 => x"00000000",
		1168 => x"00000000",
		1169 => x"00000000",
		1170 => x"00000000",
		1171 => x"00000000",
		1172 => x"00000000",
		1173 => x"00000000",
		1174 => x"00000000",
		1175 => x"00000000",
		1176 => x"00000000",
		1177 => x"00000000",
		1178 => x"00000000",
		1179 => x"00000000",
		1180 => x"00000000",
		1181 => x"00000000",
		1182 => x"00000000",
		1183 => x"00000000",
		1184 => x"00000000",
		1185 => x"00000000",
		1186 => x"00000000",
		1187 => x"00000000",
		1188 => x"00000000",
		1189 => x"00000000",
		1190 => x"00000000",
		1191 => x"00000000",
		1192 => x"00000000",
		1193 => x"00000000",
		1194 => x"00000000",
		1195 => x"00000000",
		1196 => x"00000000",
		1197 => x"00000000",
		1198 => x"00000000",
		1199 => x"00000000",
		1200 => x"00000000",
		1201 => x"00000000",
		1202 => x"00000000",
		1203 => x"00000000",
		1204 => x"00000000",
		1205 => x"00000000",
		1206 => x"00000000",
		1207 => x"00000000",
		1208 => x"00000000",
		1209 => x"00000000",
		1210 => x"00000000",
		1211 => x"00000000",
		1212 => x"00000000",
		1213 => x"00000000",
		1214 => x"00000000",
		1215 => x"00000000",
		1216 => x"00000000",
		1217 => x"00000000",
		1218 => x"00000000",
		1219 => x"00000000",
		1220 => x"00000000",
		1221 => x"00000000",
		1222 => x"00000000",
		1223 => x"00000000",
		1224 => x"00000000",
		1225 => x"00000000",
		1226 => x"00000000",
		1227 => x"00000000",
		1228 => x"00000000",
		1229 => x"00000000",
		1230 => x"00000000",
		1231 => x"00000000",
		1232 => x"00000000",
		1233 => x"00000000",
		1234 => x"00000000",
		1235 => x"00000000",
		1236 => x"00000000",
		1237 => x"00000000",
		1238 => x"00000000",
		1239 => x"00000000",
		1240 => x"00000000",
		1241 => x"00000000",
		1242 => x"00000000",
		1243 => x"00000000",
		1244 => x"00000000",
		1245 => x"00000000",
		1246 => x"00000000",
		1247 => x"00000000",
		1248 => x"00000000",
		1249 => x"00000000",
		1250 => x"00000000",
		1251 => x"00000000",
		1252 => x"00000000",
		1253 => x"00000000",
		1254 => x"00000000",
		1255 => x"00000000",
		1256 => x"00000000",
		1257 => x"00000000",
		1258 => x"00000000",
		1259 => x"00000000",
		1260 => x"00000000",
		1261 => x"00000000",
		1262 => x"00000000",
		1263 => x"00000000",
		1264 => x"00000000",
		1265 => x"00000000",
		1266 => x"00000000",
		1267 => x"00000000",
		1268 => x"00000000",
		1269 => x"00000000",
		1270 => x"00000000",
		1271 => x"00000000",
		1272 => x"00000000",
		1273 => x"00000000",
		1274 => x"00000000",
		1275 => x"00000000",
		1276 => x"00000000",
		1277 => x"00000000",
		1278 => x"00000000",
		1279 => x"00000000",
		1280 => x"00000000",
		1281 => x"00000000",
		1282 => x"00000000",
		1283 => x"00000000",
		1284 => x"00000000",
		1285 => x"00000000",
		1286 => x"00000000",
		1287 => x"00000000",
		1288 => x"00000000",
		1289 => x"00000000",
		1290 => x"00000000",
		1291 => x"00000000",
		1292 => x"00000000",
		1293 => x"00000000",
		1294 => x"00000000",
		1295 => x"00000000",
		1296 => x"00000000",
		1297 => x"00000000",
		1298 => x"00000000",
		1299 => x"00000000",
		1300 => x"00000000",
		1301 => x"00000000",
		1302 => x"00000000",
		1303 => x"00000000",
		1304 => x"00000000",
		1305 => x"00000000",
		1306 => x"00000000",
		1307 => x"00000000",
		1308 => x"00000000",
		1309 => x"00000000",
		1310 => x"00000000",
		1311 => x"00000000",
		1312 => x"00000000",
		1313 => x"00000000",
		1314 => x"00000000",
		1315 => x"00000000",
		1316 => x"00000000",
		1317 => x"00000000",
		1318 => x"00000000",
		1319 => x"00000000",
		1320 => x"00000000",
		1321 => x"00000000",
		1322 => x"00000000",
		1323 => x"00000000",
		1324 => x"00000000",
		1325 => x"00000000",
		1326 => x"00000000",
		1327 => x"00000000",
		1328 => x"00000000",
		1329 => x"00000000",
		1330 => x"00000000",
		1331 => x"00000000",
		1332 => x"00000000",
		1333 => x"00000000",
		1334 => x"00000000",
		1335 => x"00000000",
		1336 => x"00000000",
		1337 => x"00000000",
		1338 => x"00000000",
		1339 => x"00000000",
		1340 => x"00000000",
		1341 => x"00000000",
		1342 => x"00000000",
		1343 => x"00000000",
		1344 => x"00000000",
		1345 => x"00000000",
		1346 => x"00000000",
		1347 => x"00000000",
		1348 => x"00000000",
		1349 => x"00000000",
		1350 => x"00000000",
		1351 => x"00000000",
		1352 => x"00000000",
		1353 => x"00000000",
		1354 => x"00000000",
		1355 => x"00000000",
		1356 => x"00000000",
		1357 => x"00000000",
		1358 => x"00000000",
		1359 => x"00000000",
		1360 => x"00000000",
		1361 => x"00000000",
		1362 => x"00000000",
		1363 => x"00000000",
		1364 => x"00000000",
		1365 => x"00000000",
		1366 => x"00000000",
		1367 => x"00000000",
		-- Rest
		others => x"00000000"
	);


begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read -- 
			o_data <= mem(to_integer(unsigned(i_r_addr)));
			
		end if; 
	end process;

end architecture arch;